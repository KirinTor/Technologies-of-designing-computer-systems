architecture PLM_NOR of PLM_4 is
begin
 Y<=not (D or C or B or A)
 after td; 
end PLM_NOR;