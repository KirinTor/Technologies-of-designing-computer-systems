use CNetwork.all;
entity lsm_tb is
end lsm_tb;
architecture TB_ARCHITECTURE of lsm_tb is
 component LSM --?????????? ???????????? ? ?????????? ????????
 port(F : in BIT_VECTOR(1 downto 0);
 A : in BIT_VECTOR(3 downto 0);
 B : in BIT_VECTOR(3 downto 0);
 C0: in BIT;
 Y : out BIT_VECTOR(3 downto 0);
 C3: out BIT;
 Z : out BIT );
end component;
component RANDOM_GEN is
 generic(n:positive:=4; --??????????? ????????? ?????
 tp:time:=100 ns ; -- ?????? ??????????
 SEED:positive:=12345); -- ????????? ?????????
 port(CLK:out BIT;
 Y : out BIT_VECTOR(n-1 downto 0));
end component;
--??????????? ???????
signal F : BIT_VECTOR(1 downto 0):="00";
signal C0 : BIT:='0';
signal A,B : BIT_VECTOR(3 downto 0);
--??????????? ???????
signal Y1,Y2,Y : BIT_VECTOR(3 downto 0);
signal C31,C32,C, Z1,Z2,Z: BIT;
begin
G1: RANDOM_GEN --????????? ???????? ?
 generic map(n=>4,SEED=>1234)
 port map(CLK=>open,Y =>A);
G2: RANDOM_GEN --????????? ???????? ?
generic map(n=>4,SEED=>8765) 
port map(CLK=>open,Y =>B);
UUT1 :entity LSM(STR_LUT) --??????????? ??????
 port map (F => F,A => A,B => B, C0 => C0,
 Y => Y1, C3 => C31, Z => Z1);
UUT2 :entity LSM(BEH) --????????? ??????
 port map (F => F,A => A,B => B,C0 => C0,
 Y => Y2, C3 => C32, Z => Z2);
 COMP_Y: Y<=Y1 xor Y2; --??????????? ??? ????????? ???????????
 COMP_C: C<=C31 xor C32;
 COMP_Z: Z<=Z1 xor Z2;
end TB_ARCHITECTURE; 