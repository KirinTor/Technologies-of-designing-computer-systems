architecture STR_PLM of LSM is
signal c,x,yi: BIT_VECTOR(4 downto 0); --?????????? ???????
component PLM_4 is --???????????? ?????????
 --? ??????? ?????????????
 generic(td:time:=1 ns);
 port(a, b, c, d: in BIT;
 Y : out BIT);
end component;
begin
 c(0)<=C0; --??????? ???????
-- 4 ??????? LSM ---------------------------------------------------
LSM_STR:for i in 0 to 3 generate
 LNI:entity PLM_4(PLMI) port map -- ???? LNI
 (a=>A(i),b=>B(i),c=> F(0),d =>F(1), Y =>X(i));
 LNO: entity PLM_4(PLMO) port map -- ???? LNO
 (a=>C(i),b=>X(i),c=> F(0),d =>F(1), Y =>yi(i));
 LNC:entity PLM_4(PLMS) port map -- ???? LNC
 (a=>A(i),b=>B(i),c=> c(i),d =>F(0), Y =>c(i+1));
end generate;
UZ:entity PLM_4(PLM_NOR) port map(yi(3),yi(2),yi(1),yi(0),Z); --??????? ???-??
 Y<=yi(3 downto 0); -- ?????????
 C3<=c(4);
end STR_PLM; 